`define PageMask 43:28
`define VPN2 27:9
`define G 8
`define ASID 7:0
`define PFN1 49:30
`define C1 29:27
`define D1 26
`define V1 25
`define PFN0 24:5
`define C0 4:2
`define D0 1
`define V0 0
