module SRAM(
	input wire clk,  // main clock
	input wire rst,  // synchronous reset

	// SRAM interfaces
	output reg [2:0]sram_ce_n,
	output reg [2:0]sram_oe_n,
	output reg [2:0]sram_we_n,
	output reg [2:0]sram_ub_n,
	output reg [2:0]sram_lb_n,
	output reg [19:0] sram_addr,
	inout wire [47:0] sram_data,
	
	// WishBone Bus
	input wire wb_stb,  // chip select
	input wire [31:0] wb_addr,  // address
	input wire [3:0] wb_we,
	input wire [31:0] wb_din,
	output reg [31:0] wb_dout,
	output reg wb_nak
	);
	
	reg [47:0] sram_dout;
	wire [47:0] sram_din;
	assign
            sram_data = (&sram_we_n) ? {48{1'bz}} : sram_dout,
            sram_din = sram_data;
            
	localparam
		S_IDLE = 0,  // idle
		//S_START = 1,  // set address and read operation
		S_READ = 2,  // read data
		S_WRITE = 3,  // write data
		S_READ_D1 = 4,
		S_WRITE_D1 = 5;
	
	reg [2:0] state = 0;
	reg [2:0] next_state;
	reg [3:0] bus_we;
	reg [31:0] bus_din;
	
	always @(*) begin
		next_state = 0;
		case (state)
			S_IDLE: begin
				if (wb_stb)
				    if (|wb_we)
				       next_state = S_WRITE;
				    else
					   next_state = S_READ;
				else
					next_state = S_IDLE;
			end
			S_READ: begin
					next_state = S_READ_D1;
			end
			S_READ_D1: begin
			     if (wb_stb)
			        if (|wb_we)
			           next_state = S_WRITE;
			        else
			           next_state = S_READ;
			     else
			        next_state = S_IDLE;
			end
			S_WRITE: begin
                next_state = S_WRITE_D1;
            end
			S_WRITE_D1: begin
                 if (wb_stb)
                    if (|wb_we)
                       next_state = S_WRITE;
                    else
                       next_state = S_READ;
                 else
                    next_state = S_IDLE;
            end
		endcase
	end
	
	always @(posedge clk) begin
		if (rst) begin
			state <= 0;
		end
		else begin
			state <= next_state;
		end
	end
	
	always @(posedge clk) begin
		wb_nak <= 1'b1;
		sram_ce_n <= 3'b111;
		sram_oe_n <= 3'b111;
		sram_we_n <= 3'b111;
		sram_ub_n <= 3'b111;
		sram_lb_n <= 3'b111;
		sram_addr <= 20'b0;
		sram_dout <= 48'b0;
		wb_dout <= 32'b0;
		if (~rst) case (next_state)
			S_IDLE: begin
                wb_nak <= 1'b1;
			end
			S_READ: begin
			     wb_nak <= 1'b1;
			     sram_ce_n <= 3'b100;
			     sram_oe_n <= 3'b100;
			     sram_ub_n <= 3'b100;
			     sram_lb_n <= 3'b100;
			     sram_addr <= wb_addr[21:2];
			end
			S_READ_D1: begin
                wb_nak <= 1'b0;
                sram_ce_n <= sram_ce_n;
                sram_oe_n <= sram_oe_n;
                sram_ub_n <= sram_ub_n;
                sram_lb_n <= sram_lb_n;
                sram_addr <= sram_addr;
                wb_dout <= sram_din;
            end
			S_WRITE: begin
			    wb_nak <= 1'b1;
				sram_ce_n <= 3'b0;
				sram_addr <= wb_addr[21:2];
				sram_dout <= {16'b0, wb_din};
				sram_we_n <= {1'b1, ~(wb_we[3] | wb_we[2]), ~(wb_we[1] | wb_we[0])};
				sram_ub_n <= {1'b1, ~wb_we[3], ~wb_we[1]};
				sram_lb_n <= {1'b1, ~wb_we[2], ~wb_we[0]};
			end
			S_WRITE_D1: begin
			     wb_nak <= 1'b0;
			     sram_ce_n <= sram_ce_n;
			     sram_addr <= sram_addr;
			     sram_dout <= sram_dout;
			     sram_we_n <= sram_we_n;
			     sram_ub_n <= sram_ub_n;
			     sram_lb_n <= sram_lb_n;
			end
		endcase
	end
	
endmodule
